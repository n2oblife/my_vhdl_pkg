-------------------------------------------------------------------------------------------------
-- Company : ...
-- Author : nooblife
-- Licensing : MIT
-------------------------------------------------------------------------------------------------
-- Version : V1
-- Version history :
-- V1 : dd-mm-yyyy : nooblife: Creation
-------------------------------------------------------------------------------------------------
-- File name : new_file_template.vhd
-- File Creation date : dd-mm-yyyy
-- Project name : My VHDL package
-------------------------------------------------------------------------------------------------
-- Softwares :  current OS - Editor (VSCode + ...)
-------------------------------------------------------------------------------------------------
-- Description: ...
--
-- Limitations : ...
--
-------------------------------------------------------------------------------------------------
-- Naming conventions:
--
-- i_Port: Input entity port
-- o_Port: Output entity port
-- b_Port: Bidirectional entity port
-- g_My_Generic: Generic entity port
--
-- c_My_Constant: Constant definition
-- t_My_Type: Custom type definition
--
-- sc_My_Signal : Signal between components
-- My_Signal_n: Active low signal
-- v_My_Variable: Variable
-- sm_My_Signal: FSM signal
-- pkg_Param: Element Param coming from a package
--
-- My_Signal_re: Rising edge detection of My_Signal
-- My_Signal_fe: Falling edge detection of My_Signal
-- My_Signal_rX: X times registered My_Signal signal
--
-- P_Process_Name: Process
--
-------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


-------------------------------------------------------------------------------------------------
------------------------------------------ DECLARATION ------------------------------------------
-------------------------------------------------------------------------------------------------
package package_name is
-- Declaration of
    -- types and subtypes
    -- subprograms
    -- constants, signals etc.

-------------------------------------------------------------------------------------------------


-------------------------------------------------------------------------------------------------
end package_name;
-------------------------------------------------------------------------------------------------



-------------------------------------------------------------------------------------------------
--------------------------------------------- BODY ----------------------------------------------
-------------------------------------------------------------------------------------------------
package body package_name is
-- Definition of previously declared
    -- constants
    -- subprograms
-- Declaration/definition of additional
    -- types and subtypes
    -- subprograms
    -- constants, signals and shared variables

-------------------------------------------------------------------------------------------------




-------------------------------------------------------------------------------------------------
end package_name;
-------------------------------------------------------------------------------------------------